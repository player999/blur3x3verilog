library verilog;
use verilog.vl_types.all;
entity filter_tb is
end filter_tb;
